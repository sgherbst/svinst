`define MODULE_NAME mod_name_from_inc_sv
