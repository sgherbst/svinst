module A;
endmodule

modul B;
endmodule

module C;
    A I0 ();
    B I1 ();
endmodule

module D;
    X I0 ();
    Y I1 ();
endmodule
