interface b;
endinterface

module A;
endmodule

interface c;
endinterface

module E;
    c c_i ();
endmodule

interface d;
endinterface
